`ifndef _urng_vh_
`define _urng_vh_

`define URNG_BX 16

`endif //_urng_vh_
